`define DMEM_AWIDTH 18
`define NUM_BANKS 14

`include "axi_consts.vh"

`define DEBUG


//`define SOCKET_S
`define NO_AXIS

`define RAM_READ_LATENCY 5

`define MEMORY_UNIT_LATENCY 3

// MMIO addresses

`define MMIO_AW 12

`define SOCKET_MMIO_REG_SPACE 16
// These need to match software/memory_map.h
`define MMIO_KERNEL_CTRL     32'h8000_0000

`define MMIO_LSU0_CSR               32'h8000_0100
`define MMIO_LSU0_RAM_START_IDX     32'h8000_0104
`define MMIO_LSU0_RAM_BLOCK_FACTOR  32'h8000_0108
`define MMIO_LSU0_RAM_CYCLIC_FACTOR 32'h8000_010c
`define MMIO_LSU0_RAM_STRIDE        32'h8000_0110
`define MMIO_LSU0_RAM_SEG_STRIDE    32'h8000_0114
`define MMIO_LSU0_RAM_ADDR_OFFSET   32'h8000_0118
`define MMIO_LSU0_M_OFFSET_LO       32'h8000_011c
`define MMIO_LSU0_M_OFFSET_HI       32'h8000_0120
`define MMIO_LSU0_SEG_STRIDE        32'h8000_0124
`define MMIO_LSU0_SEG_COUNT         32'h8000_0128
`define MMIO_LSU0_LEN               32'h8000_012c
`define MMIO_LSU0_MODE              32'h8000_0130

`define MMIO_LSU1_CSR               32'h8000_0200
`define MMIO_LSU1_RAM_START_IDX     32'h8000_0204
`define MMIO_LSU1_RAM_BLOCK_FACTOR  32'h8000_0208
`define MMIO_LSU1_RAM_CYCLIC_FACTOR 32'h8000_020c
`define MMIO_LSU1_RAM_STRIDE        32'h8000_0210
`define MMIO_LSU1_RAM_SEG_STRIDE    32'h8000_0214
`define MMIO_LSU1_RAM_ADDR_OFFSET   32'h8000_0218
`define MMIO_LSU1_M_OFFSET_LO       32'h8000_021c
`define MMIO_LSU1_M_OFFSET_HI       32'h8000_0220
`define MMIO_LSU1_SEG_STRIDE        32'h8000_0224
`define MMIO_LSU1_SEG_COUNT         32'h8000_0228
`define MMIO_LSU1_LEN               32'h8000_022c
`define MMIO_LSU1_MODE              32'h8000_0230

`define MMIO_COMM0_MODE             32'h8000_0234
`define MMIO_COMM1_MODE             32'h8000_0238

`define MMIO_TQ_WDATA               32'h8000_0240
`define MMIO_TQ_EMPTY_N             32'h8000_0244
`define MMIO_TQ_FULL_N              32'h8000_0248

`define MMIO_CL_CFG_ENQ             32'h8000_024c

//`define MMIO_DMA0_CTRL       32'h8000_0100
//`define MMIO_DMA0_STATUS     32'h8000_0104
//`define MMIO_DMA0_IADDR_LO   32'h8000_0108
//`define MMIO_DMA0_IADDR_HI   32'h8000_010c
//`define MMIO_DMA0_EADDR_LO   32'h8000_0110
//`define MMIO_DMA0_EADDR_HI   32'h8000_0114
//`define MMIO_DMA0_LEN        32'h8000_0118
//`define MMIO_DMA0_STRIDE     32'h8000_011c
//`define MMIO_DMA0_OFFSET     32'h8000_0120
//`define MMIO_DMA0_SEG_STRIDE 32'h8000_0124
//`define MMIO_DMA0_SEG_COUNT  32'h8000_0128
//`define MMIO_DMA0_WVAL       32'h8000_0130
//`define MMIO_DMA0_MODE       32'h8000_0134
//
//`define MMIO_DMA1_CTRL       32'h8000_0200
//`define MMIO_DMA1_STATUS     32'h8000_0204
//`define MMIO_DMA1_IADDR_LO   32'h8000_0208
//`define MMIO_DMA1_IADDR_HI   32'h8000_020c
//`define MMIO_DMA1_EADDR_LO   32'h8000_0210
//`define MMIO_DMA1_EADDR_HI   32'h8000_0214
//`define MMIO_DMA1_LEN        32'h8000_0218
//`define MMIO_DMA1_STRIDE     32'h8000_021c
//`define MMIO_DMA1_OFFSET     32'h8000_0220
//`define MMIO_DMA1_SEG_STRIDE 32'h8000_0224
//`define MMIO_DMA1_SEG_COUNT  32'h8000_0228
//`define MMIO_DMA1_WVAL       32'h8000_0230
//`define MMIO_DMA1_MODE       32'h8000_0234
//
//`define MMIO_DDR_INIT_EN 32'h8000_0140

`define MMIO_SYNC(x)  (32'h8000_0150 + (x << 2))

`define MMIO_SYNC0  32'h8000_0150
`define MMIO_SYNC1  32'h8000_0154
`define MMIO_SYNC2  32'h8000_0158
`define MMIO_SYNC3  32'h8000_015c
`define MMIO_SYNC4  32'h8000_0160
`define MMIO_SYNC5  32'h8000_0164
`define MMIO_SYNC6  32'h8000_0168
`define MMIO_SYNC7  32'h8000_016c
`define MMIO_SYNC8  32'h8000_0170
`define MMIO_SYNC9  32'h8000_0174
`define MMIO_SYNC10 32'h8000_0178
`define MMIO_SYNC11 32'h8000_017c
`define MMIO_SYNC12 32'h8000_0180
`define MMIO_SYNC13 32'h8000_0184
`define MMIO_SYNC14 32'h8000_0188
`define MMIO_SYNC15 32'h8000_018c

`define MMIO_SQUEUE            32'h8000_0190
`define MMIO_SQUEUE_FULL       32'h8000_0194
`define MMIO_SQUEUE_SYNC_EMPTY 32'h8000_0198

`define MMIO_MAC_A 32'h8000_0300
`define MMIO_MAC_X 32'h8000_0304
`define MMIO_MAC_B 32'h8000_0308
`define MMIO_MAC_Y 32'h8000_030c
`define MMIO_MAC_O 32'h8000_0310

`define MMIO_MEM_UNIT_CTRL  32'h8000_0314 // {we, en}
`define MMIO_MEM_UNIT_ADDR  32'h8000_0318
`define MMIO_MEM_UNIT_WDATA 32'h8000_031c
`define MMIO_MEM_UNIT_RDATA 32'h8000_0320

`define MMIO_TASK_EMPTY 32'h8000_0344
`define MMIO_TASK_END   32'h8000_0348
`define MMIO_TASK_ADV   32'h8000_034c

`define MMIO_CPU_STATUS 32'h8000_0350

`define MMIO_CTRL_MAXI_READ             32'h8000_0354
`define MMIO_CTRL_MAXI_WRITE            32'h8000_0358
`define MMIO_CTRL_MAXI_RDATA            32'h8000_035c
`define MMIO_CTRL_MAXI_WDATA            32'h8000_0360
`define MMIO_CTRL_MAXI_SOCKET_OFFSET_LO 32'h8000_0364
`define MMIO_CTRL_MAXI_SOCKET_OFFSET_HI 32'h8000_0368

`define MMIO_SOCKET_INBOX 32'h8000_036c

`define MMIO_DMA0_WRITE_IDLE 32'h8000_0370
`define MMIO_DMA1_WRITE_IDLE 32'h8000_0374

//`define SOCKET_BASE(x)  (64'h20100000000 + 64'h40000000 * x)
`define SOCKET_BASE(x)  (64'h40000000 * (x + 1))

